LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;


ENTITY DivFreq IS
	PORT (	fin : IN STD_LOGIC; 
		fout: OUT STD_LOGIC);
END DivFreq;