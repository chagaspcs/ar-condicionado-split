LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;


ENTITY On_Off IS
	PORT (	bt : in STD_LOGIC;
		led_online : out STD_LOGIC);
END On_Off;